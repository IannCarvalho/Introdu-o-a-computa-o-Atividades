CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
34 91 1332 708
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
60 C:\Users\carva\AppData\Local\Temp\Rar$EXa0.153\CM60S\BOM.DAT
0 7
34 91 1332 708
143654930 0
0
6 Title:
5 Name:
0
0
0
31
13 Logic Switch~
5 444 390 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 443 347 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 442 302 0 1 11
0 6
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 444 262 0 1 11
0 7
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 442 143 0 1 11
0 15
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 442 96 0 1 11
0 16
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7734 0 0
0
0
13 Logic Switch~
5 130 317 0 1 11
0 20
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9914 0 0
0
0
13 Logic Switch~
5 129 272 0 1 11
0 21
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3747 0 0
0
0
13 Logic Switch~
5 132 137 0 1 11
0 26
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 C
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3549 0 0
0
0
13 Logic Switch~
5 134 96 0 1 11
0 27
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 B
-4 -29 3 -21
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7931 0 0
0
0
13 Logic Switch~
5 134 171 0 1 11
0 25
0
0 0 21360 0
2 0V
-8 -16 6 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9325 0 0
0
0
14 Logic Display~
6 808 312 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8903 0 0
0
0
5 4071~
219 732 332 0 3 22
0 4 3 2
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U3D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 -703434374
65 0 0 0 4 4 3 0
1 U
3834 0 0
0
0
5 4030~
219 639 433 0 3 22
0 6 5 3
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U7A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 -636325514
65 0 0 0 4 1 7 0
1 U
3363 0 0
0
0
5 4071~
219 636 260 0 3 22
0 7 8 4
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U3C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 -787320451
65 0 0 0 4 3 3 0
1 U
7668 0 0
0
0
5 4049~
219 501 326 0 2 22
0 6 9
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 1 6 0
1 U
4718 0 0
0
0
5 4081~
219 554 335 0 3 22
0 9 10 8
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 -636325514
65 0 0 0 4 1 5 0
1 U
3874 0 0
0
0
5 7405~
219 514 261 0 2 22
0 7 13
0
0 0 624 0
6 74LS05
-21 -24 21 -16
3 U1D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 4 1 0
1 U
6671 0 0
0
0
5 4071~
219 616 373 0 3 22
0 12 5 11
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 -552439437
65 0 0 0 4 2 3 0
1 U
3789 0 0
0
0
9 2-In AND~
219 571 270 0 3 22
0 13 6 12
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 -787320451
65 0 0 0 4 3 2 0
1 U
4871 0 0
0
0
5 4011~
219 518 115 0 3 22
0 16 15 14
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 -787320451
65 0 0 0 4 1 4 0
1 U
3750 0 0
0
0
14 Logic Display~
6 663 359 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8778 0 0
0
0
14 Logic Display~
6 589 99 0 1 2
10 14
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
538 0 0
0
0
14 Logic Display~
6 306 274 0 1 2
10 17
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6843 0 0
0
0
9 2-In AND~
219 262 294 0 3 22
0 19 18 17
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 -636325514
65 0 0 0 4 2 2 0
1 U
3136 0 0
0
0
5 7405~
219 180 317 0 2 22
0 20 18
0
0 0 624 0
6 74LS05
-21 -24 21 -16
3 U1C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 3 1 0
1 U
5950 0 0
0
0
5 7405~
219 181 272 0 2 22
0 21 19
0
0 0 624 0
6 74LS05
-21 -24 21 -16
3 U1B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 2 1 0
1 U
5670 0 0
0
0
5 4071~
219 274 112 0 3 22
0 24 23 22
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 -787320451
65 0 0 0 4 1 3 0
1 U
6828 0 0
0
0
9 2-In AND~
219 225 134 0 3 22
0 26 25 23
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 -636325514
65 0 0 0 4 1 2 0
1 U
6735 0 0
0
0
5 7405~
219 216 86 0 2 22
0 27 24
0
0 0 624 0
6 74LS05
-21 -24 21 -16
3 U1A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 1 0
1 U
8365 0 0
0
0
14 Logic Display~
6 324 99 0 1 2
22 22
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-6 -23 8 -15
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4132 0 0
0
0
30
3 1 2 0 0 4224 0 13 12 0 0 5
765 332
796 332
796 338
808 338
808 330
3 2 3 0 0 8320 0 14 13 0 0 4
672 433
711 433
711 341
719 341
3 1 4 0 0 8320 0 15 13 0 0 4
669 260
711 260
711 323
719 323
1 2 5 0 0 4224 0 1 14 0 0 4
456 390
599 390
599 442
623 442
0 1 6 0 0 8320 0 0 14 8 0 3
463 326
463 424
623 424
1 1 7 0 0 8336 0 4 15 0 0 5
456 262
456 236
615 236
615 251
623 251
3 2 8 0 0 8320 0 17 15 0 0 4
575 335
615 335
615 269
623 269
1 1 6 0 0 0 0 16 3 0 0 4
486 326
463 326
463 302
454 302
2 1 9 0 0 4224 0 16 17 0 0 2
522 326
530 326
1 2 10 0 0 4224 0 2 17 0 0 4
455 347
522 347
522 344
530 344
3 1 11 0 0 4224 0 19 22 0 0 3
649 373
663 373
663 377
1 2 5 0 0 0 0 1 19 0 0 4
456 390
595 390
595 382
603 382
3 1 12 0 0 8320 0 20 19 0 0 4
592 270
595 270
595 364
603 364
1 2 6 0 0 0 0 3 20 0 0 4
454 302
516 302
516 279
547 279
1 1 7 0 0 0 0 4 18 0 0 3
456 262
499 262
499 261
2 1 13 0 0 12416 0 18 20 0 0 4
535 261
525 261
525 261
547 261
3 1 14 0 0 4224 0 21 23 0 0 5
545 115
577 115
577 125
589 125
589 117
1 2 15 0 0 4224 0 5 21 0 0 4
454 143
486 143
486 124
494 124
1 1 16 0 0 4224 0 6 21 0 0 4
454 96
486 96
486 106
494 106
3 1 17 0 0 4224 0 25 24 0 0 3
283 294
306 294
306 292
2 2 18 0 0 4224 0 26 25 0 0 4
201 317
231 317
231 303
238 303
2 1 19 0 0 4224 0 27 25 0 0 4
202 272
231 272
231 285
238 285
1 1 20 0 0 4224 0 7 26 0 0 2
142 317
165 317
1 1 21 0 0 4224 0 8 27 0 0 2
141 272
166 272
3 1 22 0 0 4224 0 28 31 0 0 3
307 112
324 112
324 117
3 2 23 0 0 8320 0 29 28 0 0 4
246 134
252 134
252 121
261 121
2 1 24 0 0 8320 0 30 28 0 0 4
237 86
252 86
252 103
261 103
1 2 25 0 0 4224 0 11 29 0 0 4
146 171
184 171
184 143
201 143
1 1 26 0 0 4224 0 9 29 0 0 4
144 137
184 137
184 125
201 125
1 1 27 0 0 4224 0 10 30 0 0 4
146 96
187 96
187 86
201 86
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
423 203 519 227
433 211 521 227
11 Quest�o 10:
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
421 40 509 64
431 48 511 64
10 Quest�o 9:
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
107 208 195 232
117 216 197 232
10 Quest�o 8:
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
108 38 196 62
118 46 198 62
10 Quest�o 6:
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
