CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
34 91 1332 708
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
60 C:\Users\carva\AppData\Local\Temp\Rar$EXa0.601\CM60S\BOM.DAT
0 7
34 91 1332 708
143654930 0
0
6 Title:
5 Name:
0
0
0
30
13 Logic Switch~
5 569 452 0 1 11
0 13
0
0 0 21360 90
2 0V
11 0 25 8
2 V8
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 528 453 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V7
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 485 454 0 1 11
0 15
0
0 0 21360 90
2 0V
11 0 25 8
2 V6
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 49 287 0 1 11
0 17
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 50 250 0 1 11
0 18
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 50 216 0 1 11
0 19
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7734 0 0
0
0
13 Logic Switch~
5 48 107 0 1 11
0 21
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9914 0 0
0
0
13 Logic Switch~
5 49 66 0 1 11
0 22
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3747 0 0
0
0
7 Ground~
168 1215 49 0 1 3
0 2
0
0 0 53360 512
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3549 0 0
0
0
8 3-In OR~
219 1047 263 0 4 22
0 4 5 6 3
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U8A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 8 0
1 U
7931 0 0
0
0
8 2-In OR~
219 1045 332 0 3 22
0 5 6 7
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 7 0
1 U
9325 0 0
0
0
9 CC 7-Seg~
183 1178 166 0 17 19
10 3 7 5 4 3 3 3 3 2
1 0 0 1 1 1 1 1
0
0 0 21088 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 0 1 0 0 0
4 DISP
8903 0 0
0
0
7 Ground~
168 942 415 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3834 0 0
0
0
8 2-In OR~
219 817 267 0 3 22
0 9 8 5
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 681122552
65 0 0 0 4 1 7 0
1 U
3363 0 0
0
0
9 2-In AND~
219 825 178 0 3 22
0 11 10 4
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0
65 0 0 0 4 3 3 0
1 U
7668 0 0
0
0
13 2-In NAND:DM~
219 714 142 0 3 22
0 12 13 11
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U6A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 681122552
65 0 0 0 4 1 6 0
1 U
4718 0 0
0
0
9 Inverter~
13 642 312 0 2 22
0 12 14
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 2 5 0
1 U
3874 0 0
0
0
9 Inverter~
13 642 222 0 2 22
0 15 10
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 5 0
1 U
6671 0 0
0
0
9 3-In AND~
219 725 231 0 4 22
0 10 12 13 9
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 4 0
1 U
3789 0 0
0
0
9 2-In AND~
219 725 304 0 3 22
0 15 14 8
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0
65 0 0 0 4 2 3 0
1 U
4871 0 0
0
0
9 2-In AND~
219 823 375 0 3 22
0 15 12 6
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 748165885
65 0 0 0 4 1 3 0
1 U
3750 0 0
0
0
7 Ground~
168 245 245 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8778 0 0
0
0
10 3-In NAND~
219 156 236 0 4 22
0 19 18 17 16
0
0 0 624 0
6 74LS10
-21 -28 21 -20
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 2 0
1 U
538 0 0
0
0
7 Ground~
168 228 93 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6843 0 0
0
0
9 2-In XOR~
219 128 85 0 3 22
0 22 21 20
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 1771765995
65 0 0 0 4 1 1 0
1 U
3136 0 0
0
0
5 Lamp~
206 893 362 0 2 3
10 6 2
0
0 0 608 0
3 100
-10 -24 11 -16
2 L5
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
5950 0 0
0
0
5 Lamp~
206 893 254 0 2 3
11 5 2
0
0 0 608 0
3 100
-10 -24 11 -16
2 L4
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
5670 0 0
0
0
5 Lamp~
206 884 165 0 2 3
12 4 2
0
0 0 608 0
3 100
-10 -24 11 -16
2 L3
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
6828 0 0
0
0
5 Lamp~
206 217 223 0 2 3
11 16 2
0
0 0 608 0
3 100
-10 -24 11 -16
2 L1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
6735 0 0
0
0
5 Lamp~
206 194 72 0 2 3
11 20 2
0
0 0 608 0
3 100
-10 -24 11 -16
2 L2
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
8365 0 0
0
0
45
0 7 3 0 0 4096 0 0 12 2 0 3
1187 210
1187 202
1193 202
0 6 3 0 0 4096 0 0 12 3 0 4
1181 263
1181 210
1187 210
1187 202
0 5 3 0 0 8192 0 0 12 4 0 3
1157 263
1181 263
1181 202
1 4 3 0 0 8320 0 12 10 0 0 3
1157 202
1157 263
1080 263
8 0 3 0 0 0 0 12 0 0 6 2
1199 202
1199 202
5 6 3 0 0 0 0 12 12 0 0 4
1181 202
1222 202
1222 202
1187 202
1 9 2 0 0 12288 0 9 12 0 0 6
1215 43
1215 39
1229 39
1229 115
1178 115
1178 124
4 0 4 0 0 8192 0 12 0 0 14 4
1175 202
1175 217
1021 217
1021 222
0 3 5 0 0 12432 0 0 12 11 0 6
1012 264
992 264
992 210
1168 210
1168 202
1169 202
0 2 6 0 0 4096 0 0 11 12 0 3
1006 272
1006 341
1032 341
0 1 5 0 0 0 0 0 11 13 0 3
1013 264
1013 323
1032 323
0 3 6 0 0 8320 0 0 10 21 0 3
875 375
875 272
1034 272
0 2 5 0 0 128 0 0 10 20 0 4
877 267
877 264
1035 264
1035 263
0 1 4 0 0 8320 0 0 10 19 0 5
863 178
863 222
1022 222
1022 254
1034 254
2 3 7 0 0 4224 0 12 11 0 0 3
1163 202
1163 332
1078 332
0 1 2 0 0 0 0 0 13 18 0 2
942 374
942 409
2 0 2 0 0 8192 0 28 0 0 18 4
896 178
943 178
943 267
942 267
2 2 2 0 0 8320 0 27 26 0 0 6
905 267
942 267
942 374
913 374
913 375
905 375
3 1 4 0 0 0 0 15 28 0 0 2
846 178
872 178
3 1 5 0 0 0 0 14 27 0 0 2
850 267
881 267
3 1 6 0 0 0 0 21 26 0 0 2
844 375
881 375
3 2 8 0 0 4224 0 20 14 0 0 4
746 304
796 304
796 276
804 276
4 1 9 0 0 4224 0 19 14 0 0 4
746 231
796 231
796 258
804 258
0 2 10 0 0 8320 0 0 15 33 0 3
680 222
680 187
801 187
3 1 11 0 0 4224 0 16 15 0 0 4
747 142
783 142
783 169
801 169
0 1 12 0 0 8192 0 0 16 32 0 3
529 231
529 133
695 133
0 2 13 0 0 8192 0 0 16 31 0 3
570 245
570 151
695 151
2 2 14 0 0 4224 0 17 20 0 0 4
663 312
693 312
693 313
701 313
0 1 12 0 0 0 0 0 17 32 0 2
529 312
627 312
0 1 15 0 0 4096 0 0 20 34 0 2
486 295
701 295
1 3 13 0 0 4224 0 1 19 0 0 3
570 439
570 240
701 240
0 2 12 0 0 8192 0 0 19 36 0 3
529 394
529 231
701 231
2 1 10 0 0 0 0 18 19 0 0 2
663 222
701 222
0 1 15 0 0 0 0 0 18 35 0 3
486 376
486 222
627 222
1 1 15 0 0 8320 0 3 21 0 0 3
486 441
486 366
799 366
1 2 12 0 0 8320 0 2 21 0 0 3
529 440
529 384
799 384
2 1 2 0 0 0 0 29 22 0 0 3
229 236
245 236
245 239
4 1 16 0 0 4224 0 23 29 0 0 2
183 236
205 236
1 3 17 0 0 8320 0 4 23 0 0 5
61 287
61 268
124 268
124 245
132 245
1 2 18 0 0 8320 0 5 23 0 0 3
62 250
62 236
132 236
1 1 19 0 0 4224 0 6 23 0 0 4
62 216
124 216
124 227
132 227
2 1 2 0 0 0 0 30 24 0 0 5
206 85
215 85
215 79
228 79
228 87
3 1 20 0 0 4224 0 25 30 0 0 2
161 85
182 85
1 2 21 0 0 4224 0 7 25 0 0 4
60 107
107 107
107 94
112 94
1 1 22 0 0 4224 0 8 25 0 0 4
61 66
107 66
107 76
112 76
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
